library verilog;
use verilog.vl_types.all;
entity Multiplicadores_vlg_vec_tst is
end Multiplicadores_vlg_vec_tst;

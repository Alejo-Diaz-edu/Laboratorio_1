library verilog;
use verilog.vl_types.all;
entity pruebacontador_vlg_check_tst is
    port(
        Cout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end pruebacontador_vlg_check_tst;

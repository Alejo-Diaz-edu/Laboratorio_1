library verilog;
use verilog.vl_types.all;
entity pruebacontador is
    port(
        Cout            : out    vl_logic;
        clock           : in     vl_logic
    );
end pruebacontador;

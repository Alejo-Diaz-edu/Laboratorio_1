-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Oct 30 14:55:48 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY I2E_Maquina_De_Estado IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        fin_dir : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        SDA : IN STD_LOGIC := '0';
        Hab_Dir : OUT STD_LOGIC;
        Hab_Dat : OUT STD_LOGIC;
        ACK : OUT STD_LOGIC
    );
END I2E_Maquina_De_Estado;

ARCHITECTURE BEHAVIOR OF I2E_Maquina_De_Estado IS
    TYPE type_fstate IS (RoW,ACK_State,Guarda_Dat,Guarda_dir,Idle);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,fin_dir,soy,fin_dato,SDA)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Idle;
            Hab_Dir <= '0';
            Hab_Dat <= '0';
            ACK <= '0';
        ELSE
            Hab_Dir <= '0';
            Hab_Dat <= '0';
            ACK <= '0';
            CASE fstate IS
                WHEN RoW =>
                    reg_fstate <= ACK_State;

                    Hab_Dir <= '0';
                    Hab_Dir <= '0';
                    Hab_Dir <= '0';
                WHEN ACK_State =>
                    reg_fstate <= Guarda_Dat;

                    Hab_Dat <= '0';

                    ACK <= '1';

                    Hab_Dir <= '0';
                WHEN Guarda_Dat =>
                    IF ((fin_dato = '1')) THEN
                        reg_fstate <= Idle;
                    ELSIF ((fin_dato = '0')) THEN
                        reg_fstate <= Guarda_Dat;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_Dat;
                    END IF;

                    Hab_Dat <= '1';

                    ACK <= '0';

                    Hab_Dir <= '0';
                WHEN Guarda_dir =>
                    IF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= RoW;
                    ELSIF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Idle;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guarda_dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_dir;
                    END IF;

                    Hab_Dat <= '0';

                    ACK <= '0';

                    Hab_Dir <= '1';
                WHEN Idle =>
                    IF ((SDA = '0')) THEN
                        reg_fstate <= Guarda_dir;
                    ELSIF ((SDA = '1')) THEN
                        reg_fstate <= Idle;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Idle;
                    END IF;

                    Hab_Dat <= '0';

                    ACK <= '0';

                    Hab_Dir <= '0';
                WHEN OTHERS => 
                    Hab_Dir <= 'X';
                    Hab_Dat <= 'X';
                    ACK <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;

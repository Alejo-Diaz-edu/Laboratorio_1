library verilog;
use verilog.vl_types.all;
entity MultiplicadorSS_vlg_vec_tst is
end MultiplicadorSS_vlg_vec_tst;

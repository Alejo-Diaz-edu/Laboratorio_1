library verilog;
use verilog.vl_types.all;
entity MultiplicadorSS_vlg_check_tst is
    port(
        R0              : in     vl_logic;
        R1              : in     vl_logic;
        R2              : in     vl_logic;
        R3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MultiplicadorSS_vlg_check_tst;

-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Thu Oct 23 16:37:22 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY MultiplicadorCS IS 
	PORT
	(
		B0 :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		R0 :  OUT  STD_LOGIC;
		R1 :  OUT  STD_LOGIC;
		R2 :  OUT  STD_LOGIC;
		R3 :  OUT  STD_LOGIC;
		SIGNO :  OUT  STD_LOGIC
	);
END MultiplicadorCS;

ARCHITECTURE bdf_type OF MultiplicadorCS IS 

COMPONENT fulladder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 Cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_45 <= '1';
SYNTHESIZED_WIRE_48 <= '0';
SYNTHESIZED_WIRE_8 <= '0';
SYNTHESIZED_WIRE_17 <= '1';
SYNTHESIZED_WIRE_21 <= '0';
SYNTHESIZED_WIRE_25 <= '1';
SYNTHESIZED_WIRE_51 <= '1';
SYNTHESIZED_WIRE_52 <= '1';



SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_44;


PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	R0 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	R0 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	R0 <= SYNTHESIZED_WIRE_1;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_49 <= SYNTHESIZED_WIRE_46 AND SYNTHESIZED_WIRE_44;


b2v_inst17 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_47,
		 B => SYNTHESIZED_WIRE_48,
		 Cin => SYNTHESIZED_WIRE_5,
		 S => SYNTHESIZED_WIRE_19,
		 Cout => SYNTHESIZED_WIRE_22);


b2v_inst18 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_6,
		 B => SYNTHESIZED_WIRE_49,
		 Cin => SYNTHESIZED_WIRE_8,
		 S => SYNTHESIZED_WIRE_38,
		 Cout => SYNTHESIZED_WIRE_11);


b2v_inst19 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_9,
		 B => SYNTHESIZED_WIRE_49,
		 Cin => SYNTHESIZED_WIRE_11,
		 S => SYNTHESIZED_WIRE_41,
		 Cout => SYNTHESIZED_WIRE_14);


b2v_inst20 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_12,
		 B => SYNTHESIZED_WIRE_49,
		 Cin => SYNTHESIZED_WIRE_14,
		 S => SYNTHESIZED_WIRE_36);


b2v_inst21 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_15,
		 B => SYNTHESIZED_WIRE_48,
		 Cin => SYNTHESIZED_WIRE_17,
		 S => SYNTHESIZED_WIRE_18,
		 Cout => SYNTHESIZED_WIRE_5);




SYNTHESIZED_WIRE_15 <= NOT(SYNTHESIZED_WIRE_43);



SYNTHESIZED_WIRE_47 <= NOT(SYNTHESIZED_WIRE_46);



SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_18 AND SYNTHESIZED_WIRE_50;


SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_50;


b2v_inst28 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_47,
		 B => SYNTHESIZED_WIRE_21,
		 Cin => SYNTHESIZED_WIRE_22,
		 S => SYNTHESIZED_WIRE_23);



SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_46 XOR SYNTHESIZED_WIRE_50;



SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_50;


PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_25)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '0';
ELSIF (SYNTHESIZED_WIRE_25 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_43 <= A0;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_46 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_46 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_46 <= A1;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_44 <= B0;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_51)
BEGIN
IF (SYNTHESIZED_WIRE_51 = '0') THEN
	SYNTHESIZED_WIRE_50 <= '0';
ELSIF (SYNTHESIZED_WIRE_51 = '0') THEN
	SYNTHESIZED_WIRE_50 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_50 <= B1;
END IF;
END PROCESS;





PROCESS(CLK,SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_52 = '0') THEN
	SIGNO <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	SIGNO <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SIGNO <= SYNTHESIZED_WIRE_33;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_52 = '0') THEN
	R3 <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	R3 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	R3 <= SYNTHESIZED_WIRE_36;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_52 = '0') THEN
	R1 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	R1 <= SYNTHESIZED_WIRE_38;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_52 = '0') THEN
	R2 <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	R2 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	R2 <= SYNTHESIZED_WIRE_41;
END IF;
END PROCESS;



END bdf_type;
library verilog;
use verilog.vl_types.all;
entity pruebacontador_vlg_vec_tst is
end pruebacontador_vlg_vec_tst;

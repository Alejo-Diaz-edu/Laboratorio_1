library verilog;
use verilog.vl_types.all;
entity I2E_completo_vlg_vec_tst is
end I2E_completo_vlg_vec_tst;
